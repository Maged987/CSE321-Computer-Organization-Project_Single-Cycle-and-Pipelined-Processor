
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.records_pkg.all;
use work.segm_mips_const_pkg.all;

entity WRITE_BACK is
port( 
	--Entradas
	RESET			: in STD_LOGIC;					--Reset
	WB			    : in WB_CTRL_REG;				
	READ_DATA		: in STD_LOGIC_VECTOR (INST_SIZE-1 downto 0);	-- data that comes from data memory
	ADDRESS			: in STD_LOGIC_VECTOR (INST_SIZE-1 downto 0);	-- data that comes from ALU
	WRITE_REG		: in STD_LOGIC_VECTOR (ADDR_SIZE-1 downto 0);	--from control unit to register files		
	
	RegWrite		: out STD_LOGIC;				
	WRITE_REG_OUT	: out STD_LOGIC_VECTOR (ADDR_SIZE-1 downto 0);	--Register destination address
	WRITE_DATA		: out STD_LOGIC_VECTOR (INST_SIZE-1 downto 0)	--Data to write into register file
);
end WRITE_BACK;

architecture WRITE_BACK_ARC of WRITE_BACK is 
begin

	MUX_WB: 
		process(RESET,WB.RegWrite,WRITE_REG,WB.MemtoReg,ADDRESS,READ_DATA)
		begin
			if( RESET = '1') then
				RegWrite <= '0';
				WRITE_REG_OUT <= "00000"; 
				WRITE_DATA <= ZERO32b; 
			else
				RegWrite <= WB.RegWrite;
				WRITE_REG_OUT <= WRITE_REG;
			 	if( WB.MemtoReg = '0') then
			 		WRITE_DATA <= ADDRESS; 
			 	else
			 		WRITE_DATA <= READ_DATA;
			 	end if;
			end if;
		 end process MUX_WB;
		 
end WRITE_BACK_ARC;
